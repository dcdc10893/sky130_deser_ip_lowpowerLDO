** sch_path: /home/dcdc/xschem-src/Work1/chipalooza2024/sky130_deser_ip_lowpowerLDO_upload/cace/test_temp4.sch
**.subckt test_temp4
Vref Vref VSUB DC {VVref}
Vena Vena VSUB DC {VVena}
Vvss vss VSUB DC {Vvss}
Rout out VSUB {Rout} m=1
Cout out VSUB {Cout} m=1
Vvdd vdd VSUB DC {Vvdd}
RSUB VSUB GND 0.01 m=1
x1 Vref out vdd vss vss VSUB Vena sky130_deser_ip_lowpowerLDO
**** begin user architecture code

.control
op
ac dec 20 1 1e6
let vog = 20 * log(V(out))+40
meas vres MAX vog
echo $&vres > {simpath}/{filename}_{N}.data

setplot new
plot db(V(out))+40

quit
.endc



* CACE gensim simulation file {filename}_{N}
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the amplifier under condition of static input


.lib {PDK_ROOT}/{PDK}/libs.tech/combined/sky130.lib.spice {corner}

.option TEMP={temperature}
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1


**** end user architecture code
**.ends

* expanding   symbol:  xschem/sky130_deser_ip_lowpowerLDO.sym # of pins=7
** sym_path: /home/dcdc/xschem-src/Work1/chipalooza2024/sky130_deser_ip_lowpowerLDO_upload/xschem/sky130_deser_ip_lowpowerLDO.sym
** sch_path: /home/dcdc/xschem-src/Work1/chipalooza2024/sky130_deser_ip_lowpowerLDO_upload/xschem/sky130_deser_ip_lowpowerLDO.sch
.subckt sky130_deser_ip_lowpowerLDO Vref Vout avdd dvdd avss dvss ena
*.ipin avdd
*.ipin dvss
*.ipin dvdd
*.ipin avss
*.ipin ena
*.ipin Vref
*.opin Vout
XR10 Vfed Vout avdd sky130_fd_pr__res_xhigh_po_5p73 L=5.73*150 mult=1 m=1
XR4 avss Vfed avdd sky130_fd_pr__res_xhigh_po_5p73 L=5.73*300 mult=1 m=1
XR8 avss net3 avdd sky130_fd_pr__res_xhigh_po_5p73 L=5.73*500 mult=1 m=1
XC4 Vout_fb3 net4 sky130_fd_pr__cap_mim_m3_2 W=10 L=20 MF=1 m=1
R9 net4 Vout_fb1 sky130_fd_pr__res_generic_l1 W=1 L=19 m=1
XM6 net3 net3 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5*1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)
+ * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net1 net3 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)
+ * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vout_fb1 net3 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)
+ * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 Vout_fb3 Vfed net1 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=14 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf
+ * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 Vref net1 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=14 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)
+ * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 Vout Vout_fb1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=80 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf
+ * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM8 Vout_fb3 net2 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=13 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf
+ * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 Vout_fb1 Vout_fb3 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf
+ * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 net2 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=13 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)
+ * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 Vout_fb2 ena Vout_fb1 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2.7*1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)
+ * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 Vout_fb2 ena dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1*1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf
+ * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R2 avss dvss sky130_fd_pr__res_generic_l1 W=3 L=1 m=1
.ends

.GLOBAL GND
.end
